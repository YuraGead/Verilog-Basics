// радуга на семисегменте буквой

module lab
(
input [2:0] sw,
output [6:0] segm
);

assign segm = (sw == 3'b001) ? ~7'b1110111 : 
				 ((sw == 3'b010) ? ~7'b0111111 :
				 ((sw == 3'b011) ? ~7'b1101110 :
				 ((sw == 3'b100) ? ~7'b1111101 :
				 ((sw == 3'b101) ? ~7'b1111111 :
				 ((sw == 3'b110) ? ~7'b0000110 :
				 ((sw == 3'b111) ? ~7'b0111110 :
				 ~7'b0000000))))));

				 
				 
//0 = 0
//1 = ~7'b1110111 /R
//2 = ~7'b0111111 /O
//3 = ~7'b1101110 /Y
//4 = ~7'b1111101 /G
//5 = ~7'b1111111 /B
//6 = ~7'b0000110 /I
//7 = ~7'b0111110 /V
endmodule 